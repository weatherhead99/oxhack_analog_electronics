* /home/danw/Documents/oxhack_analog_electronics/schematics/VCO/VCO.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon 20 Nov 2017 23:14:27 GMT

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0
.include 2N7000.REV0.SP3
.include TL081.301
.param control_v =3

* Sheet Name: /
XU1  16 17 1 3 13 TL081		;Node Sequence Spec.<3,2,7,4,6>
C2  1 14 10nF		
C3  3 14 10nF		
XU2  15 13 1 3 5 TL081		;Node Sequence Spec.<3,2,7,4,6>
C4  1 14 10nF		
C5  3 14 10nF		
R1  16 4 100k		
R2  16 14 49.9k		
R3  17 4 100k		
C1  13 17 10nF		
XQ1  14 5 12 2n7000		
R4  17 12 49.9k		
R6  15 14 100k		
R7  5 15 100k		
R5  1 15 380k		
V1  1 14 +12		
V2  2 3 +12		
V3  4 14 control_v		

.end
